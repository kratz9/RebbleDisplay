`timescale 1 ns / 1 ps

module rebble_screen
  (
   input  wire  reset,
   input  wire  cs,
   output wire  miso
   input  wire  mosi,
   input  wire  sck,
	 
   output wire reset_done,
   output wire intn
   );
   
   






  endmodule
